//*****************************************************************
// Name:    <Your Name> 
// Date:    <Term Year>
// File     function04.v
// Purp:    f04 logic function
//
// Assisted by: Christopher Coulston Spring 2020
//
// Academic Integrity Statement: I certify that, while others may have
// assisted me in brain storming, debugging and validating this program,
// the program itself is my own work. I understand that submitting code
// which is the work of other individuals is a violation of the course
// Academic Integrity Policy and may result in a zero credit for the
// assignment, course failure and a report to the Academic Dishonesty
// Board. I also understand that if I knowingly give my original work to
// another individual that it could also result in a zero credit for the
// assignment, course failure and a report to the Academic Dishonesty
// Board.
//*****************************************************************
module function04(a, b, c, f04);

    input  a, b, c;
    output f04;

    // Wires are signals that begin and end inside the module
    wire o1, a1, a2;

    // Complete the following lines of verilog code

    assign o1 =
    assign a1 =
    assign a2 =
    assign f04 =

endmodule
