//------------------------------------------
//	Name:	Chris Coulston
// Date:	Spring 2020
// File:	sevent_segment
//	Purp:	Hex to 7-segment converter
//------------------------------------------
//
//		Active low LEDs on segments
//
//				 hex[0]
//				 -----
//	hex[5]	|		|	hex[1]
//				|		|	
//				 -----	hex[6]
//	hex[4]	|		|
//				|		|	hex[2]
//				 -----
//				 hex[3]
//
//------------------------------------------

module sevenSegment(X, S);
	output reg [6:0] S;
	input wire [3:0] X;
	
	always @(*)
		case (X)
			4'b0000: S = 7'b1000000;	// 0 = 1000000
			4'b0001: S = 7'b1111001;   // 1 = 1111001
			4'b0010: S = 7'b0100100;   // 2 = 0100100
			4'b0011: S = 7'b0110000;   // 3 = 0110000
			4'b0100: S = 7'b0011001;   // 4 = 0011001
			4'b0101: S = 7'b0010010;   // 5 = 0010010
			4'b0110: S = 7'b0000010;   // 6 = 0000010
			4'b0111: S = 7'b1111000;   // 7 = 1111000
			4'b1000: S = 7'b0000000;   // 8 = 0000000
			4'b1001: S = 7'b0011000;   // 9 = 0011000
			4'b1010: S = 7'b0001000;   // A = 0001000
			4'b1011: S = 7'b0000011;   // b = 0000011
			4'b1100: S = 7'b1000110;   // C = 1000110
			4'b1101: S = 7'b0100001;   // d = 0100001
			4'b1110: S = 7'b0000110;   // E = 0000110
			4'b1111: S = 7'b0001110;   // F = 0001110
		endcase
endmodule
