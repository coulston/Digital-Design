//*****************************************************************
// Name:     
// Date:     
// Lab:     03
// Purp:    playToSeven
//
// Assisted: The entire EENG 284 class
// Assisted by: Dr. Christopher Coulston
//------------------------------------------------
//
//	Active low LEDs on segments
//
//            seg[0]
//		        ------
//	  seg[5]  |      |   seg[1]
//           |      |	
//            ------ seg[6]
//   seg[4]  |      |
//           |      |   seg[2]
//            ------
//            seg[3]
//
//------------------------------------------
module playToSeven (pPlay, sevenSeg);



endmodule
