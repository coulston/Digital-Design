//*****************************************************************
// Name:    <Your Name>
// Date:    <Term Year>
// File:    lfsrStart.c
// Purp:    lfsr module
//
// Assisted: Christopher Coulston and Thomas MacDougall Spring 2023
//
// Academic Integrity Statement: I certify that, while others may have
// assisted me in brain storming, debugging and validating this program,
// the program itself is my own work. I understand that submitting code
// which is the work of other individuals is a violation of the course
// Academic Integrity Policy and may result in a zero credit for the
// assignment, course failure and a report to the Academic Dishonesty
// Board. I also understand that if I knowingly give my original work to
// another individual that it could also result in a zero credit for the
// assignment, course failure and a report to the Academic Dishonesty
// Board.
//*****************************************************************
module lfsr(inputSeed, outputRand);

    // Put variable decelaration here

    assign outputRand[0] =
    assign outputRand[1] =
    assign outputRand[2] =
    assign outputRand[3] =

endmodule
