//*****************************************************************
// Name:    <Your Name>
// Date:    
// Lab:     03
// Purp:    winLoose
//
// Assisted: The entire EENG 284 class
// Assisted by: Dr. Christopher Coulston
//------------------------------------------------
//
//	Active low LEDs on segments
//
//            seg[0]
//		        ------
//	  seg[5]  |      |   seg[1]
//           |      |	
//            ------ seg[6]
//   seg[4]  |      |
//           |      |   seg[2]
//            ------
//            seg[3]
//
//
//	button nominally logic 1, when pressed equals 0
//
//*****************************************************************
module winLose(p1Play, p2Play, playButton, sevenSeg);







endmodule
