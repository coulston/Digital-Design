//*****************************************************************
// Name:    <Your Name>
// Date:    Spring 2020
// Lab:     03
// Purp:    winLoose
//
// Assisted: The entire EENG 383 class
// Assisted by: Dr. Vibhuti Dave
//
// Academic Integrity Statement: I certify that, while others may have
// assisted me in brain storming, debugging and validating this program,
// the program itself is my own work. I understand that submitting code
// which is the work of other individuals is a violation of the course
// Academic Integrity Policy and may result in a zero credit for the
// assignment, course failure and a report to the Academic Dishonesty
// Board. I also understand that if I knowingly give my original work to
// another individual that it could also result in a zero credit for the
// assignment, course failure and a report to the Academic Dishonesty
// Board.
//
//------------------------------------------
//
//	Active low LEDs on segments
//
//            seg[0]
//		        ------
//	  seg[5]  |      |   seg[1]
//           |      |
//            ------ seg[6]
//   seg[4]  |      |
//           |      |   seg[2]
//            ------
//            seg[3]
//
//
//	button nominally logic 1, when pressed equals 0
//
//*****************************************************************
module winLose(p1Play, p2Play, playButton, sevenSeg);







endmodule
