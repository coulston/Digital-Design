//*****************************************************************
// Name:    <Your Name>
// Date:     
// Lab:     03
// Purp:    rpsGame
//
// Assisted: The entire EENG 284 class
// Assisted by: Dr. Christopher Coulston
//------------------------------------------------
//*****************************************************************
module rpsGame(p1Throw, p1SevenSeg, p2Throw, p2SevenSeg, playButton, winLoseSeg);
	

	     
    onesToDense p1o2d(p1Throw, p1Dense);


endmodule
