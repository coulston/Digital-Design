//*****************************************************************
// Name:    <Your Name> 
// Date:    <Term Year>
// File:    function02.v
// Purp:    Realize f02 = a’ + bc’
//
// Assisted by: Christopher Coulston Spring 2020
//
// Academic Integrity Statement: I certify that, while others may have
// assisted me in brain storming, debugging and validating this program,
// the program itself is my own work. I understand that submitting code
// which is the work of other individuals is a violation of the course
// Academic Integrity Policy and may result in a zero credit for the
// assignment, course failure and a report to the Academic Dishonesty
// Board. I also understand that if I knowingly give my original work to
// another individual that it could also result in a zero credit for the
// assignment, course failure and a report to the Academic Dishonesty
// Board.
//*****************************************************************
module function02 (a, b, c, f02);

    input  a, b, c;
    output f02;

    // Complete the following line of verilog code
    // Use the logic operators and parenthesis

    assign f02 =

endmodule
