//*****************************************************************
// Name:     
// Date:     
// Lab:     03
// Purp:    playToSeven
//
// Assisted: The entire EENG 284 class
// Assisted by: Dr. Christopher Coulston
//------------------------------------------------
//    play[1] = 
//    play[0] = 
//*****************************************************************
module onesToDense (throw, play);




endmodule
